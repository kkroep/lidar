LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY gfz2lino IS
    PORT(
        SIGNAL GFZ_LP       : IN std_logic_vector(1 TO 70);
        SIGNAL GFZ_LN       : IN std_logic_vector(1 TO 70);
        SIGNAL GFZ_RP       : IN std_logic_vector(1 TO 70);
        SIGNAL GFZ_RN       : IN std_logic_vector(1 TO 70);
        
        SIGNAL LINO_MAIN    : OUT std_logic_vector(255 DOWNTO 0);
        SIGNAL LINO_AUX     : OUT std_logic_vector(7 DOWNTO 0)
    );
END ENTITY gfz2lino;

ARCHITECTURE arch OF gfz2lino IS
    SIGNAL aux : std_logic_vector(8 DOWNTO 1);
    SIGNAL o : std_logic_vector(256 DOWNTO 1);
BEGIN
    LINO_AUX <= aux;
    LINO_MAIN <= o;

    --Pixel input wiring
    aux(1) <= GFZ_RN(66);
    aux(2) <= GFZ_RN(68);
    aux(3) <= GFZ_RN(45);
    aux(4) <= GFZ_RN(44);
    aux(5) <= GFZ_LP(70);
    aux(6) <= GFZ_LP(69);
    aux(7) <= GFZ_LN(41);
    aux(8) <= GFZ_LP(48);

    o(1) <= GFZ_RN(69);
    o(2) <= GFZ_LN(65);
    o(3) <= GFZ_RN(61);
    o(4) <= GFZ_LN(64);
    o(5) <= GFZ_RN(67);
    o(6) <= GFZ_LN(63);
    o(7) <= GFZ_RN(62);
    o(8) <= GFZ_LP(66);
    o(9) <= GFZ_RN(70);
    o(10) <= GFZ_LP(62);
    o(11) <= GFZ_RP(64);
    o(12) <= GFZ_LP(68);
    o(13) <= GFZ_RP(62);
    o(14) <= GFZ_LN(62);
    o(15) <= GFZ_RN(65);
    o(16) <= GFZ_LP(67);
    o(17) <= GFZ_RP(67);
    o(18) <= GFZ_LN(61);
    o(19) <= GFZ_RN(63);
    o(20) <= GFZ_LP(61);
    o(21) <= GFZ_RP(63);
    o(22) <= GFZ_LP(40);
    o(23) <= GFZ_RP(61);
    o(24) <= GFZ_LN(69);
    o(25) <= GFZ_RP(68);
    o(26) <= GFZ_LP(65);
    o(27) <= GFZ_RN(64);
    o(28) <= GFZ_LP(63);
    o(29) <= GFZ_RP(65);
    o(30) <= GFZ_LP(64);
    o(31) <= GFZ_RN(36);
    o(32) <= GFZ_LN(33);
    o(33) <= GFZ_RN(38);
    o(34) <= GFZ_LN(39);
    o(35) <= GFZ_RP(36);
    o(36) <= GFZ_LN(30);
    o(37) <= GFZ_RP(39);
    o(38) <= GFZ_LP(39);
    o(39) <= GFZ_RP(35);
    o(40) <= GFZ_LP(29);
    o(41) <= GFZ_RP(30);
    o(42) <= GFZ_LN(40);
    o(43) <= GFZ_RP(26);
    o(44) <= GFZ_LP(28);
    o(45) <= GFZ_RN(28);
    o(46) <= GFZ_LN(32);
    o(47) <= GFZ_RP(34);
    o(48) <= GFZ_LP(27);
    o(49) <= GFZ_RP(21);
    o(50) <= GFZ_LN(31);
    o(51) <= GFZ_RP(32);
    o(52) <= GFZ_LN(25);
    o(53) <= GFZ_RN(21);
    o(54) <= GFZ_LN(35);
    o(55) <= GFZ_RP(33);
    o(56) <= GFZ_LN(24);
    o(57) <= GFZ_RN(22);
    o(58) <= GFZ_LP(31);
    o(59) <= GFZ_RP(31);
    o(60) <= GFZ_LN(23);
    o(61) <= GFZ_RP(25);
    o(62) <= GFZ_LP(37);
    o(63) <= GFZ_RN(39);
    o(64) <= GFZ_LP(23);
    o(65) <= GFZ_RN(25);
    o(66) <= GFZ_LP(38);
    o(67) <= GFZ_RN(37);
    o(68) <= GFZ_LP(22);
    o(69) <= GFZ_RP(23);
    o(70) <= GFZ_LN(37);
    o(71) <= GFZ_RP(27);
    o(72) <= GFZ_LN(21);
    o(73) <= GFZ_RP(16);
    o(74) <= GFZ_LN(26);
    o(75) <= GFZ_RN(20);
    o(76) <= GFZ_LP(21);
    o(77) <= GFZ_RN(24);
    o(78) <= GFZ_LP(30);
    o(79) <= GFZ_RN(17);
    o(80) <= GFZ_LN(20);
    o(81) <= GFZ_RP(20);
    o(82) <= GFZ_LN(17);
    o(83) <= GFZ_RN(16);
    o(84) <= GFZ_LP(24);
    o(85) <= GFZ_RN(23);
    o(86) <= GFZ_LN(19);
    o(87) <= GFZ_RN(33);
    o(88) <= GFZ_LN(18);
    o(89) <= GFZ_RP(18);
    o(90) <= GFZ_LN(22);
    o(91) <= GFZ_RP(37);
    o(92) <= GFZ_LN(68);
    o(93) <= GFZ_RP(69);
    o(94) <= GFZ_LN(36);
    o(95) <= GFZ_RN(40);
    o(96) <= GFZ_LN(29);
    o(97) <= GFZ_RP(38);
    o(98) <= GFZ_LN(38);
    o(99) <= GFZ_RP(40);
    o(100) <= GFZ_LN(27);
    o(101) <= GFZ_RP(29);
    o(102) <= GFZ_LP(36);
    o(103) <= GFZ_RN(32);
    o(104) <= GFZ_LN(28);
    o(105) <= GFZ_RP(28);
    o(106) <= GFZ_LP(34);
    o(107) <= GFZ_RN(35);
    o(108) <= GFZ_LN(67);
    o(109) <= GFZ_RP(70);
    o(110) <= GFZ_LP(35);
    o(111) <= GFZ_RN(31);
    o(112) <= GFZ_LP(26);
    o(113) <= GFZ_RP(22);
    o(114) <= GFZ_LN(34);
    o(115) <= GFZ_RN(34);
    o(116) <= GFZ_LP(25);
    o(117) <= GFZ_RP(24);
    o(118) <= GFZ_LP(33);
    o(119) <= GFZ_RN(27);
    o(120) <= GFZ_LN(16);
    o(121) <= GFZ_RP(17);
    o(122) <= GFZ_LN(9);
    o(123) <= GFZ_RN(30);
    o(124) <= GFZ_LN(66);
    o(125) <= GFZ_RP(66);
    o(126) <= GFZ_LP(32);
    o(127) <= GFZ_RN(26);
    o(128) <= GFZ_LP(19);
    o(129) <= GFZ_RP(19);
    o(130) <= GFZ_LP(6);
    o(131) <= GFZ_RN(8);
    o(132) <= GFZ_LN(50);
    o(133) <= GFZ_RN(47);
    o(134) <= GFZ_LP(8);
    o(135) <= GFZ_RN(29);
    o(136) <= GFZ_LN(12);
    o(137) <= GFZ_RP(11);
    o(138) <= GFZ_LP(7);
    o(139) <= GFZ_RN(1);
    o(140) <= GFZ_LP(14);
    o(141) <= GFZ_RP(13);
    o(142) <= GFZ_LN(4);
    o(143) <= GFZ_RN(5);
    o(144) <= GFZ_LN(7);
    o(145) <= GFZ_RP(9);
    o(146) <= GFZ_LP(1);
    o(147) <= GFZ_RN(4);
    o(148) <= GFZ_LN(49);
    o(149) <= GFZ_RN(50);
    o(150) <= GFZ_LP(3);
    o(151) <= GFZ_RN(2);
    o(152) <= GFZ_LP(10);
    o(153) <= GFZ_RP(8);
    o(154) <= GFZ_LP(2);
    o(155) <= GFZ_RN(3);
    o(156) <= GFZ_LP(9);
    o(157) <= GFZ_RP(1);
    o(158) <= GFZ_LN(60);
    o(159) <= GFZ_RN(57);
    o(160) <= GFZ_LP(60);
    o(161) <= GFZ_RP(5);
    o(162) <= GFZ_LP(57);
    o(163) <= GFZ_RN(60);
    o(164) <= GFZ_LN(46);
    o(165) <= GFZ_RN(49);
    o(166) <= GFZ_LP(20);
    o(167) <= GFZ_RP(7);
    o(168) <= GFZ_LN(5);
    o(169) <= GFZ_RP(15);
    o(170) <= GFZ_LN(15);
    o(171) <= GFZ_RN(19);
    o(172) <= GFZ_LP(16);
    o(173) <= GFZ_RP(14);
    o(174) <= GFZ_LN(13);
    o(175) <= GFZ_RP(12);
    o(176) <= GFZ_LP(17);
    o(177) <= GFZ_RN(18);
    o(178) <= GFZ_LN(14);
    o(179) <= GFZ_RN(9);
    o(180) <= GFZ_LP(18);
    o(181) <= GFZ_RN(11);
    o(182) <= GFZ_LN(11);
    o(183) <= GFZ_RP(2);
    o(184) <= GFZ_LN(2);
    o(185) <= GFZ_RP(6);
    o(186) <= GFZ_LP(15);
    o(187) <= GFZ_RP(52);
    o(188) <= GFZ_LP(55);
    o(189) <= GFZ_RN(12);
    o(190) <= GFZ_LP(13);
    o(191) <= GFZ_RP(58);
    o(192) <= GFZ_LN(53);
    o(193) <= GFZ_RN(15);
    o(194) <= GFZ_LN(8);
    o(195) <= GFZ_RP(51);
    o(196) <= GFZ_LN(56);
    o(197) <= GFZ_RP(10);
    o(198) <= GFZ_LP(12);
    o(199) <= GFZ_RP(3);
    o(200) <= GFZ_LP(5);
    o(201) <= GFZ_RN(14);
    o(202) <= GFZ_LP(11);
    o(203) <= GFZ_RP(59);
    o(204) <= GFZ_LN(57);
    o(205) <= GFZ_RN(13);
    o(206) <= GFZ_LN(6);
    o(207) <= GFZ_RP(60);
    o(208) <= GFZ_LP(4);
    o(209) <= GFZ_RN(6);
    o(210) <= GFZ_LN(10);
    o(211) <= GFZ_RP(57);
    o(212) <= GFZ_LN(1);
    o(213) <= GFZ_RN(7);
    o(214) <= GFZ_LN(3);
    o(215) <= GFZ_RP(55);
    o(216) <= GFZ_LN(58);
    o(217) <= GFZ_RN(10);
    o(218) <= GFZ_LN(59);
    o(219) <= GFZ_RN(56);
    o(220) <= GFZ_LP(59);
    o(221) <= GFZ_RP(4);
    o(222) <= GFZ_LP(58);
    o(223) <= GFZ_RN(59);
    o(224) <= GFZ_LN(52);
    o(225) <= GFZ_RP(56);
    o(226) <= GFZ_LP(56);
    o(227) <= GFZ_RN(51);
    o(228) <= GFZ_LP(54);
    o(229) <= GFZ_RP(54);
    o(230) <= GFZ_LN(51);
    o(231) <= GFZ_RN(52);
    o(232) <= GFZ_LP(47);
    o(233) <= GFZ_RN(48);
    o(234) <= GFZ_LN(55);
    o(235) <= GFZ_RN(58);
    o(236) <= GFZ_LN(48);
    o(237) <= GFZ_RP(53);
    o(238) <= GFZ_LN(54);
    o(239) <= GFZ_RN(55);
    o(240) <= GFZ_LP(49);
    o(241) <= GFZ_RP(49);
    o(242) <= GFZ_LP(53);
    o(243) <= GFZ_RN(54);
    o(244) <= GFZ_LN(47);
    o(245) <= GFZ_RP(50);
    o(246) <= GFZ_LP(51);
    o(247) <= GFZ_RP(46);
    o(248) <= GFZ_LN(42);
    o(249) <= GFZ_RP(48);
    o(250) <= GFZ_LP(50);
    o(251) <= GFZ_RN(53);
    o(252) <= GFZ_LP(46);
    o(253) <= GFZ_RP(47);
    o(254) <= GFZ_LP(52);
    o(255) <= GFZ_RN(46);
    o(256) <= GFZ_LN(43);
END ARCHITECTURE arch;
        